module tb_flanger();

// Your testbench goes here.

endmodule: tb_flanger

// Any other simulation-only modules you need

