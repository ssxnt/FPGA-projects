`timescale 1ps / 1ps

module tb_syn_task1();

    

endmodule: tb_syn_task1
