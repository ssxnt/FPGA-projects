module tb_rtl_init();

// Your testbench goes here.

endmodule: tb_rtl_init
