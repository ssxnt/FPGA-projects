module tb_music();

// Your testbench goes here.

endmodule: tb_music

// Any other simulation-only modules you need

