module tb_syn_crack();

// Your testbench goes here.

endmodule: tb_syn_crack
