module tb_syn_task2();

// Your testbench goes here.

endmodule: tb_syn_task2
