module tb_rtl_arc4();

// Your testbench goes here.

endmodule: tb_rtl_arc4
