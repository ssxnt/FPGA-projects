module tb_rtl_task2();

// Your testbench goes here.

endmodule: tb_rtl_task2
