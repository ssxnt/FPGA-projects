module tb_rtl_ksa();

// Your testbench goes here.

endmodule: tb_rtl_ksa
