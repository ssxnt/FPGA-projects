module tb_rtl_doublecrack();

// Your testbench goes here.

endmodule: tb_rtl_doublecrack
