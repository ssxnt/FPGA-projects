module tb_syn_doublecrack();

// Your testbench goes here.

endmodule: tb_syn_doublecrack
