module tb_syn_ksa();

// Your testbench goes here.

endmodule: tb_syn_ksa
