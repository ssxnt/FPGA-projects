module tb_syn_task4();

// Your testbench goes here.

endmodule: tb_syn_task4
