    Mac OS X            	   2   �      �                                      ATTR       �   �   (                  �     com.apple.lastuseddate#PS       �     com.apple.quarantine yVe    �M�5    q/0081;65075623;Chrome; 