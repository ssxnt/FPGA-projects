module tb_rtl_prga();

// Your testbench goes here.

endmodule: tb_rtl_prga
