    Mac OS X            	   2   ~      �                                      ATTR       �   �                     �     com.apple.quarantine q/0081;65075623;Chrome; 