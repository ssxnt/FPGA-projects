module tb_rtl_task1();

// Your testbench goes here.

endmodule: tb_rtl_task1
