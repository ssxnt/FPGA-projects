module tb_syn_task1();

// Your testbench goes here.

endmodule: tb_syn_task1
