module tb_syn_init();

// Your testbench goes here.

endmodule: tb_syn_init
