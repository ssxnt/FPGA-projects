module tb_rtl_task5();

// Your testbench goes here.

endmodule: tb_rtl_task5
